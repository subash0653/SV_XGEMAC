interface xgemac_rst_interface(input clk);

  logic rst;

  initial begin
    $display("XGEMAC_RST_INTERFACE");
  end

endinterface: xgemac_rst_interface
