interface xgemac_clk_interface();

  logic clk;

  initial begin
    $display("XGEMAC_CLK_INTERFACE");
  end

endinterface: xgemac_clk_interface
